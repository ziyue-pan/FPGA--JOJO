
module ROM_music(
	input clk,
	input [7:0] address,
	output reg [7:0] note
);

always @(posedge clk)
case(address)
0: note<= 8'd33;
1: note<= 8'd33;
2: note<= 8'd33;
3: note<= 8'd33;
4: note<= 8'd33;
5: note<= 8'd33;
6: note<= 8'd32;
7: note<= 8'd32;
8: note<= 8'd32;
9: note<= 8'd32;
10: note<= 8'd32;
11: note<= 8'd32;
12: note<= 8'd00;
13: note<= 8'd00;
14: note<= 8'd29;
15: note<= 8'd31;
16: note<= 8'd32;
17: note<= 8'd32;
18: note<= 8'd32;
19: note<= 8'd31;
20: note<= 8'd31;
21: note<= 8'd31;
22: note<= 8'd29;
23: note<= 8'd29;
24: note<= 8'd28;
25: note<= 8'd28;
26: note<= 8'd28;
27: note<= 8'd29;
28: note<= 8'd29;
29: note<= 8'd29;
30: note<= 8'd31;
31: note<= 8'd31;
32: note<= 8'd33;
33: note<= 8'd33;
34: note<= 8'd33;
35: note<= 8'd33;
36: note<= 8'd00;
37: note<= 8'd00;
38: note<= 8'd26;
39: note<= 8'd26;
40: note<= 8'd26;
41: note<= 8'd26;
42: note<= 8'd26;
43: note<= 8'd26;
44: note<= 8'd00;
45: note<= 8'd00;
46: note<= 8'd26;
47: note<= 8'd27;
48: note<= 8'd29;
49: note<= 8'd29;
50: note<= 8'd29;
51: note<= 8'd31;
52: note<= 8'd31;
53: note<= 8'd31;
54: note<= 8'd29;
55: note<= 8'd29;
56: note<= 8'd28;
57: note<= 8'd28;
58: note<= 8'd28;
59: note<= 8'd24;
60: note<= 8'd24;
61: note<= 8'd24;
62: note<= 8'd22;
63: note<= 8'd22;
64: note<= 8'd33;
65: note<= 8'd33;
66: note<= 8'd33;
67: note<= 8'd33;
68: note<= 8'd00;
69: note<= 8'd00;
70: note<= 8'd32;
71: note<= 8'd32;
72: note<= 8'd32;
73: note<= 8'd32;
74: note<= 8'd32;
75: note<= 8'd32;
76: note<= 8'd29;
77: note<= 8'd29;
78: note<= 8'd31;
79: note<= 8'd31;
80: note<= 8'd32;
81: note<= 8'd32;
82: note<= 8'd32;
83: note<= 8'd31;
84: note<= 8'd31;
85: note<= 8'd31;
86: note<= 8'd29;
87: note<= 8'd29;
88: note<= 8'd28;
89: note<= 8'd28;
90: note<= 8'd28;
91: note<= 8'd29;
92: note<= 8'd29;
93: note<= 8'd29;
94: note<= 8'd31;
95: note<= 8'd31;
96: note<= 8'd33;
97: note<= 8'd33;
98: note<= 8'd33;
99: note<= 8'd33;
100: note<= 8'd00;
101: note<= 8'd00;
102: note<= 8'd26;
103: note<= 8'd26;
104: note<= 8'd26;
105: note<= 8'd26;
106: note<= 8'd26;
107: note<= 8'd26;
108: note<= 8'd26;
109: note<= 8'd26;
110: note<= 8'd28;
111: note<= 8'd28;
112: note<= 8'd29;
113: note<= 8'd29;
114: note<= 8'd29;
115: note<= 8'd22;
116: note<= 8'd22;
117: note<= 8'd22;
118: note<= 8'd33;
119: note<= 8'd33;
120: note<= 8'd32;
121: note<= 8'd32;
122: note<= 8'd32;
123: note<= 8'd29;
124: note<= 8'd29;
125: note<= 8'd29;
126: note<= 8'd25;
127: note<= 8'd25;
128: note<= 8'd26;
129: note<= 8'd26;
130: note<= 8'd26;
131: note<= 8'd26;
132: note<= 8'd26;
133: note<= 8'd24;
134: note<= 8'd24;
135: note<= 8'd26;
136: note<= 8'd26;
137: note<= 8'd29;
138: note<= 8'd29;
139: note<= 8'd26;
140: note<= 8'd26;
141: note<= 8'd33;
142: note<= 8'd24;
143: note<= 8'd24;
144: note<= 8'd26;
145: note<= 8'd26;
146: note<= 8'd26;
147: note<= 8'd26;
148: note<= 8'd26;
149: note<= 8'd24;
150: note<= 8'd24;
151: note<= 8'd26;
152: note<= 8'd26;
153: note<= 8'd32;
154: note<= 8'd32;
155: note<= 8'd31;
156: note<= 8'd31;
157: note<= 8'd29;
158: note<= 8'd24;
159: note<= 8'd24;

	default: note <= 8'd0;
endcase
endmodule