module ROM_Wall(
	input clk,
	input [4:0] row,
	input [3:0] col,
	output reg [11:0] rgb
);

(* rom_style = "block" *)

//signal declaration
reg [4:0] row_reg;
reg [3:0] col_reg;

always @(posedge clk) begin
	row_reg <= row;
	col_reg <= col;
end

always @*
	case ({row_reg, col_reg})
		9'b000000000: rgb = 12'b011011011110;
		9'b000000001: rgb = 12'b000000000000;
		9'b000000010: rgb = 12'b000000000000;
		9'b000000011: rgb = 12'b000000000000;
		9'b000000100: rgb = 12'b000000000000;
		9'b000000101: rgb = 12'b000000000000;
		9'b000000110: rgb = 12'b000000000000;
		9'b000000111: rgb = 12'b000000000000;
		9'b000001000: rgb = 12'b000000000000;
		9'b000001001: rgb = 12'b000000000000;
		9'b000001010: rgb = 12'b000000000000;
		9'b000001011: rgb = 12'b000000000000;
		9'b000001100: rgb = 12'b000000000000;
		9'b000001101: rgb = 12'b000000000000;
		9'b000001110: rgb = 12'b000000000000;
		9'b000001111: rgb = 12'b011011011110;
		9'b000010000: rgb = 12'b000000000000;
		9'b000010001: rgb = 12'b000000000000;
		9'b000010010: rgb = 12'b110011001101;
		9'b000010011: rgb = 12'b110011001101;
		9'b000010100: rgb = 12'b110011001101;
		9'b000010101: rgb = 12'b110011001101;
		9'b000010110: rgb = 12'b110011001101;
		9'b000010111: rgb = 12'b110011001101;
		9'b000011000: rgb = 12'b110011001101;
		9'b000011001: rgb = 12'b110011001101;
		9'b000011010: rgb = 12'b110011001101;
		9'b000011011: rgb = 12'b110011001101;
		9'b000011100: rgb = 12'b100110011001;
		9'b000011101: rgb = 12'b100110011001;
		9'b000011110: rgb = 12'b000000000000;
		9'b000011111: rgb = 12'b000000000000;
		9'b000100000: rgb = 12'b000000000000;
		9'b000100001: rgb = 12'b000000000000;
		9'b000100010: rgb = 12'b110011001101;
		9'b000100011: rgb = 12'b110011001101;
		9'b000100100: rgb = 12'b110011001101;
		9'b000100101: rgb = 12'b110011001101;
		9'b000100110: rgb = 12'b110011001101;
		9'b000100111: rgb = 12'b110011001101;
		9'b000101000: rgb = 12'b110011001101;
		9'b000101001: rgb = 12'b100110011001;
		9'b000101010: rgb = 12'b100110011001;
		9'b000101011: rgb = 12'b100110011001;
		9'b000101100: rgb = 12'b100110011001;
		9'b000101101: rgb = 12'b100110011001;
		9'b000101110: rgb = 12'b100110011001;
		9'b000101111: rgb = 12'b000000000000;

		9'b000110000: rgb = 12'b000000000000;
		9'b000110001: rgb = 12'b110011001101;
		9'b000110010: rgb = 12'b110011001101;
		9'b000110011: rgb = 12'b110011001101;
		9'b000110100: rgb = 12'b100110011001;
		9'b000110101: rgb = 12'b100110011001;
		9'b000110110: rgb = 12'b110011001101;
		9'b000110111: rgb = 12'b110011001101;
		9'b000111000: rgb = 12'b110011001101;
		9'b000111001: rgb = 12'b100110011001;
		9'b000111010: rgb = 12'b100110011001;
		9'b000111011: rgb = 12'b100110011001;
		9'b000111100: rgb = 12'b100110011001;
		9'b000111101: rgb = 12'b100110011001;
		9'b000111110: rgb = 12'b010101010101;
		9'b000111111: rgb = 12'b000000000000;

		9'b001000000: rgb = 12'b000000000000;
		9'b001000001: rgb = 12'b110011001101;
		9'b001000010: rgb = 12'b110011001101;
		9'b001000011: rgb = 12'b110011001101;
		9'b001000100: rgb = 12'b100110011001;
		9'b001000101: rgb = 12'b100110011001;
		9'b001000110: rgb = 12'b110011001101;
		9'b001000111: rgb = 12'b110011001101;
		9'b001001000: rgb = 12'b110011001101;
		9'b001001001: rgb = 12'b100110011001;
		9'b001001010: rgb = 12'b100110011001;
		9'b001001011: rgb = 12'b100110011001;
		9'b001001100: rgb = 12'b100110011001;
		9'b001001101: rgb = 12'b100110011001;
		9'b001001110: rgb = 12'b010101010101;
		9'b001001111: rgb = 12'b000000000000;

		9'b001010000: rgb = 12'b000000000000;
		9'b001010001: rgb = 12'b110011001101;
		9'b001010010: rgb = 12'b110011001101;
		9'b001010011: rgb = 12'b100110011001;
		9'b001010100: rgb = 12'b100110011001;
		9'b001010101: rgb = 12'b100110011001;
		9'b001010110: rgb = 12'b100110011001;
		9'b001010111: rgb = 12'b100110011001;
		9'b001011000: rgb = 12'b100110011001;
		9'b001011001: rgb = 12'b100110011001;
		9'b001011010: rgb = 12'b100110011001;
		9'b001011011: rgb = 12'b100110011001;
		9'b001011100: rgb = 12'b100110011001;
		9'b001011101: rgb = 12'b100110011001;
		9'b001011110: rgb = 12'b010101010101;
		9'b001011111: rgb = 12'b000000000000;

		9'b001100000: rgb = 12'b000000000000;
		9'b001100001: rgb = 12'b110011001101;
		9'b001100010: rgb = 12'b110011001101;
		9'b001100011: rgb = 12'b100110011001;
		9'b001100100: rgb = 12'b100110011001;
		9'b001100101: rgb = 12'b100110011001;
		9'b001100110: rgb = 12'b110011001101;
		9'b001100111: rgb = 12'b110011001101;
		9'b001101000: rgb = 12'b100110011001;
		9'b001101001: rgb = 12'b100110011001;
		9'b001101010: rgb = 12'b100110011001;
		9'b001101011: rgb = 12'b100110011001;
		9'b001101100: rgb = 12'b010101010101;
		9'b001101101: rgb = 12'b010101010101;
		9'b001101110: rgb = 12'b010101010101;
		9'b001101111: rgb = 12'b000000000000;

		9'b001110000: rgb = 12'b000000000000;
		9'b001110001: rgb = 12'b110011001101;
		9'b001110010: rgb = 12'b110011001101;
		9'b001110011: rgb = 12'b100110011001;
		9'b001110100: rgb = 12'b100110011001;
		9'b001110101: rgb = 12'b100110011001;
		9'b001110110: rgb = 12'b110011001101;
		9'b001110111: rgb = 12'b110011001101;
		9'b001111000: rgb = 12'b100110011001;
		9'b001111001: rgb = 12'b100110011001;
		9'b001111010: rgb = 12'b010101010101;
		9'b001111011: rgb = 12'b010101010101;
		9'b001111100: rgb = 12'b100110011001;
		9'b001111101: rgb = 12'b010101010101;
		9'b001111110: rgb = 12'b010101010101;
		9'b001111111: rgb = 12'b000000000000;

		9'b010000000: rgb = 12'b000000000000;
		9'b010000001: rgb = 12'b100110011001;
		9'b010000010: rgb = 12'b100110011001;
		9'b010000011: rgb = 12'b100110011001;
		9'b010000100: rgb = 12'b100110011001;
		9'b010000101: rgb = 12'b100110011001;
		9'b010000110: rgb = 12'b110011001101;
		9'b010000111: rgb = 12'b110011001101;
		9'b010001000: rgb = 12'b100110011001;
		9'b010001001: rgb = 12'b100110011001;
		9'b010001010: rgb = 12'b010101010101;
		9'b010001011: rgb = 12'b010101010101;
		9'b010001100: rgb = 12'b100110011001;
		9'b010001101: rgb = 12'b010101010101;
		9'b010001110: rgb = 12'b010101010101;
		9'b010001111: rgb = 12'b000000000000;

		9'b010010000: rgb = 12'b000000000000;
		9'b010010001: rgb = 12'b100110011001;
		9'b010010010: rgb = 12'b100110011001;
		9'b010010011: rgb = 12'b010101010101;
		9'b010010100: rgb = 12'b100110011001;
		9'b010010101: rgb = 12'b100110011001;
		9'b010010110: rgb = 12'b100110011001;
		9'b010010111: rgb = 12'b100110011001;
		9'b010011000: rgb = 12'b100110011001;
		9'b010011001: rgb = 12'b100110011001;
		9'b010011010: rgb = 12'b010101010101;
		9'b010011011: rgb = 12'b010101010101;
		9'b010011100: rgb = 12'b010101010101;
		9'b010011101: rgb = 12'b010101010101;
		9'b010011110: rgb = 12'b010101010101;
		9'b010011111: rgb = 12'b000000000000;

		9'b010100000: rgb = 12'b000000000000;
		9'b010100001: rgb = 12'b100110011001;
		9'b010100010: rgb = 12'b100110011001;
		9'b010100011: rgb = 12'b100110011001;
		9'b010100100: rgb = 12'b100110011001;
		9'b010100101: rgb = 12'b100110011001;
		9'b010100110: rgb = 12'b100110011001;
		9'b010100111: rgb = 12'b100110011001;
		9'b010101000: rgb = 12'b010101010101;
		9'b010101001: rgb = 12'b010101010101;
		9'b010101010: rgb = 12'b010101010101;
		9'b010101011: rgb = 12'b010101010101;
		9'b010101100: rgb = 12'b010101010101;
		9'b010101101: rgb = 12'b010101010101;
		9'b010101110: rgb = 12'b010101010101;
		9'b010101111: rgb = 12'b000000000000;

		9'b010110000: rgb = 12'b000000000000;
		9'b010110001: rgb = 12'b100110011001;
		9'b010110010: rgb = 12'b100110011001;
		9'b010110011: rgb = 12'b010101010101;
		9'b010110100: rgb = 12'b110011001101;
		9'b010110101: rgb = 12'b110011001101;
		9'b010110110: rgb = 12'b010101010101;
		9'b010110111: rgb = 12'b010101010101;
		9'b010111000: rgb = 12'b010101010101;
		9'b010111001: rgb = 12'b010101010101;
		9'b010111010: rgb = 12'b010101010101;
		9'b010111011: rgb = 12'b100110011001;
		9'b010111100: rgb = 12'b100110011001;
		9'b010111101: rgb = 12'b010101010101;
		9'b010111110: rgb = 12'b010101010101;
		9'b010111111: rgb = 12'b000000000000;

		9'b011000000: rgb = 12'b000000000000;
		9'b011000001: rgb = 12'b010101010101;
		9'b011000010: rgb = 12'b010101010101;
		9'b011000011: rgb = 12'b010101010101;
		9'b011000100: rgb = 12'b110011001101;
		9'b011000101: rgb = 12'b110011001101;
		9'b011000110: rgb = 12'b010101010101;
		9'b011000111: rgb = 12'b010101010101;
		9'b011001000: rgb = 12'b010101010101;
		9'b011001001: rgb = 12'b010101010101;
		9'b011001010: rgb = 12'b010101010101;
		9'b011001011: rgb = 12'b100110011001;
		9'b011001100: rgb = 12'b100110011001;
		9'b011001101: rgb = 12'b010101010101;
		9'b011001110: rgb = 12'b010101010101;
		9'b011001111: rgb = 12'b000000000000;

		9'b011010000: rgb = 12'b000000000000;
		9'b011010001: rgb = 12'b010101010101;
		9'b011010010: rgb = 12'b010101010101;
		9'b011010011: rgb = 12'b010101010101;
		9'b011010100: rgb = 12'b010101010101;
		9'b011010101: rgb = 12'b010101010101;
		9'b011010110: rgb = 12'b010101010101;
		9'b011010111: rgb = 12'b010101010101;
		9'b011011000: rgb = 12'b010101010101;
		9'b011011001: rgb = 12'b010101010101;
		9'b011011010: rgb = 12'b010101010101;
		9'b011011011: rgb = 12'b010101010101;
		9'b011011100: rgb = 12'b010101010101;
		9'b011011101: rgb = 12'b010101010101;
		9'b011011110: rgb = 12'b000000000000;
		9'b011011111: rgb = 12'b000000000000;

		9'b011100000: rgb = 12'b000000000000;
		9'b011100001: rgb = 12'b000000000000;
		9'b011100010: rgb = 12'b010101010101;
		9'b011100011: rgb = 12'b010101010101;
		9'b011100100: rgb = 12'b010101010101;
		9'b011100101: rgb = 12'b010101010101;
		9'b011100110: rgb = 12'b010101010101;
		9'b011100111: rgb = 12'b010101010101;
		9'b011101000: rgb = 12'b010101010101;
		9'b011101001: rgb = 12'b010101010101;
		9'b011101010: rgb = 12'b010101010101;
		9'b011101011: rgb = 12'b010101010101;
		9'b011101100: rgb = 12'b010101010101;
		9'b011101101: rgb = 12'b000000000000;
		9'b011101110: rgb = 12'b000000000000;
		9'b011101111: rgb = 12'b000000000000;

		9'b011110000: rgb = 12'b011011011110;
		9'b011110001: rgb = 12'b000000000000;
		9'b011110010: rgb = 12'b000000000000;
		9'b011110011: rgb = 12'b000000000000;
		9'b011110100: rgb = 12'b000000000000;
		9'b011110101: rgb = 12'b000000000000;
		9'b011110110: rgb = 12'b000000000000;
		9'b011110111: rgb = 12'b000000000000;
		9'b011111000: rgb = 12'b000000000000;
		9'b011111001: rgb = 12'b000000000000;
		9'b011111010: rgb = 12'b000000000000;
		9'b011111011: rgb = 12'b000000000000;
		9'b011111100: rgb = 12'b000000000000;
		9'b011111101: rgb = 12'b000000000000;
		9'b011111110: rgb = 12'b000000000000;
		9'b011111111: rgb = 12'b011011011110;

		9'b100000000: rgb = 12'b011011011110;
		9'b100000001: rgb = 12'b000000000000;
		9'b100000010: rgb = 12'b000000000000;
		9'b100000011: rgb = 12'b000000000000;
		9'b100000100: rgb = 12'b000000000000;
		9'b100000101: rgb = 12'b000000000000;
		9'b100000110: rgb = 12'b000000000000;
		9'b100000111: rgb = 12'b000000000000;
		9'b100001000: rgb = 12'b000000000000;
		9'b100001001: rgb = 12'b000000000000;
		9'b100001010: rgb = 12'b000000000000;
		9'b100001011: rgb = 12'b000000000000;
		9'b100001100: rgb = 12'b000000000000;
		9'b100001101: rgb = 12'b000000000000;
		9'b100001110: rgb = 12'b000000000000;
		9'b100001111: rgb = 12'b011011011110;

		9'b100010000: rgb = 12'b000000000000;
		9'b100010001: rgb = 12'b000000000000;
		9'b100010010: rgb = 12'b110011001101;
		9'b100010011: rgb = 12'b110011001101;
		9'b100010100: rgb = 12'b110011001101;
		9'b100010101: rgb = 12'b110011001101;
		9'b100010110: rgb = 12'b110011001101;
		9'b100010111: rgb = 12'b110011001101;
		9'b100011000: rgb = 12'b110011001101;
		9'b100011001: rgb = 12'b110011001101;
		9'b100011010: rgb = 12'b110011001101;
		9'b100011011: rgb = 12'b110011001101;
		9'b100011100: rgb = 12'b100110011001;
		9'b100011101: rgb = 12'b100110011001;
		9'b100011110: rgb = 12'b000000000000;
		9'b100011111: rgb = 12'b000000000000;

		9'b100100000: rgb = 12'b000000000000;
		9'b100100001: rgb = 12'b000000000000;
		9'b100100010: rgb = 12'b110011001101;
		9'b100100011: rgb = 12'b110011001101;
		9'b100100100: rgb = 12'b110011001101;
		9'b100100101: rgb = 12'b110011001101;
		9'b100100110: rgb = 12'b110011001101;
		9'b100100111: rgb = 12'b110011001101;
		9'b100101000: rgb = 12'b110011001101;
		9'b100101001: rgb = 12'b100110011001;
		9'b100101010: rgb = 12'b100110011001;
		9'b100101011: rgb = 12'b100110011001;
		9'b100101100: rgb = 12'b100110011001;
		9'b100101101: rgb = 12'b100110011001;
		9'b100101110: rgb = 12'b100110011001;
		9'b100101111: rgb = 12'b000000000000;

		9'b100110000: rgb = 12'b000000000000;
		9'b100110001: rgb = 12'b110011001101;
		9'b100110010: rgb = 12'b110011001101;
		9'b100110011: rgb = 12'b110011001101;
		9'b100110100: rgb = 12'b100110011001;
		9'b100110101: rgb = 12'b100110011001;
		9'b100110110: rgb = 12'b110011001101;
		9'b100110111: rgb = 12'b110011001101;
		9'b100111000: rgb = 12'b110011001101;
		9'b100111001: rgb = 12'b100110011001;
		9'b100111010: rgb = 12'b100110011001;
		9'b100111011: rgb = 12'b100110011001;
		9'b100111100: rgb = 12'b100110011001;
		9'b100111101: rgb = 12'b100110011001;
		9'b100111110: rgb = 12'b010101010101;
		9'b100111111: rgb = 12'b000000000000;

		9'b101000000: rgb = 12'b000000000000;
		9'b101000001: rgb = 12'b110011001101;
		9'b101000010: rgb = 12'b110011001101;
		9'b101000011: rgb = 12'b110011001101;
		9'b101000100: rgb = 12'b100110011001;
		9'b101000101: rgb = 12'b100110011001;
		9'b101000110: rgb = 12'b110011001101;
		9'b101000111: rgb = 12'b110011001101;
		9'b101001000: rgb = 12'b110011001101;
		9'b101001001: rgb = 12'b100110011001;
		9'b101001010: rgb = 12'b100110011001;
		9'b101001011: rgb = 12'b100110011001;
		9'b101001100: rgb = 12'b100110011001;
		9'b101001101: rgb = 12'b100110011001;
		9'b101001110: rgb = 12'b010101010101;
		9'b101001111: rgb = 12'b000000000000;

		9'b101010000: rgb = 12'b000000000000;
		9'b101010001: rgb = 12'b110011001101;
		9'b101010010: rgb = 12'b110011001101;
		9'b101010011: rgb = 12'b100110011001;
		9'b101010100: rgb = 12'b100110011001;
		9'b101010101: rgb = 12'b100110011001;
		9'b101010110: rgb = 12'b100110011001;
		9'b101010111: rgb = 12'b100110011001;
		9'b101011000: rgb = 12'b100110011001;
		9'b101011001: rgb = 12'b100110011001;
		9'b101011010: rgb = 12'b100110011001;
		9'b101011011: rgb = 12'b100110011001;
		9'b101011100: rgb = 12'b100110011001;
		9'b101011101: rgb = 12'b100110011001;
		9'b101011110: rgb = 12'b010101010101;
		9'b101011111: rgb = 12'b000000000000;

		9'b101100000: rgb = 12'b000000000000;
		9'b101100001: rgb = 12'b110011001101;
		9'b101100010: rgb = 12'b110011001101;
		9'b101100011: rgb = 12'b100110011001;
		9'b101100100: rgb = 12'b100110011001;
		9'b101100101: rgb = 12'b100110011001;
		9'b101100110: rgb = 12'b110011001101;
		9'b101100111: rgb = 12'b110011001101;
		9'b101101000: rgb = 12'b100110011001;
		9'b101101001: rgb = 12'b100110011001;
		9'b101101010: rgb = 12'b100110011001;
		9'b101101011: rgb = 12'b100110011001;
		9'b101101100: rgb = 12'b010101010101;
		9'b101101101: rgb = 12'b010101010101;
		9'b101101110: rgb = 12'b010101010101;
		9'b101101111: rgb = 12'b000000000000;

		9'b101110000: rgb = 12'b000000000000;
		9'b101110001: rgb = 12'b110011001101;
		9'b101110010: rgb = 12'b110011001101;
		9'b101110011: rgb = 12'b100110011001;
		9'b101110100: rgb = 12'b100110011001;
		9'b101110101: rgb = 12'b100110011001;
		9'b101110110: rgb = 12'b110011001101;
		9'b101110111: rgb = 12'b110011001101;
		9'b101111000: rgb = 12'b100110011001;
		9'b101111001: rgb = 12'b100110011001;
		9'b101111010: rgb = 12'b010101010101;
		9'b101111011: rgb = 12'b010101010101;
		9'b101111100: rgb = 12'b100110011001;
		9'b101111101: rgb = 12'b010101010101;
		9'b101111110: rgb = 12'b010101010101;
		9'b101111111: rgb = 12'b000000000000;

		9'b110000000: rgb = 12'b000000000000;
		9'b110000001: rgb = 12'b100110011001;
		9'b110000010: rgb = 12'b100110011001;
		9'b110000011: rgb = 12'b100110011001;
		9'b110000100: rgb = 12'b100110011001;
		9'b110000101: rgb = 12'b100110011001;
		9'b110000110: rgb = 12'b110011001101;
		9'b110000111: rgb = 12'b110011001101;
		9'b110001000: rgb = 12'b100110011001;
		9'b110001001: rgb = 12'b100110011001;
		9'b110001010: rgb = 12'b010101010101;
		9'b110001011: rgb = 12'b010101010101;
		9'b110001100: rgb = 12'b100110011001;
		9'b110001101: rgb = 12'b010101010101;
		9'b110001110: rgb = 12'b010101010101;
		9'b110001111: rgb = 12'b000000000000;

		9'b110010000: rgb = 12'b000000000000;
		9'b110010001: rgb = 12'b100110011001;
		9'b110010010: rgb = 12'b100110011001;
		9'b110010011: rgb = 12'b010101010101;
		9'b110010100: rgb = 12'b100110011001;
		9'b110010101: rgb = 12'b100110011001;
		9'b110010110: rgb = 12'b100110011001;
		9'b110010111: rgb = 12'b100110011001;
		9'b110011000: rgb = 12'b100110011001;
		9'b110011001: rgb = 12'b100110011001;
		9'b110011010: rgb = 12'b010101010101;
		9'b110011011: rgb = 12'b010101010101;
		9'b110011100: rgb = 12'b010101010101;
		9'b110011101: rgb = 12'b010101010101;
		9'b110011110: rgb = 12'b010101010101;
		9'b110011111: rgb = 12'b000000000000;

		9'b110100000: rgb = 12'b000000000000;
		9'b110100001: rgb = 12'b100110011001;
		9'b110100010: rgb = 12'b100110011001;
		9'b110100011: rgb = 12'b100110011001;
		9'b110100100: rgb = 12'b100110011001;
		9'b110100101: rgb = 12'b100110011001;
		9'b110100110: rgb = 12'b100110011001;
		9'b110100111: rgb = 12'b100110011001;
		9'b110101000: rgb = 12'b010101010101;
		9'b110101001: rgb = 12'b010101010101;
		9'b110101010: rgb = 12'b010101010101;
		9'b110101011: rgb = 12'b010101010101;
		9'b110101100: rgb = 12'b010101010101;
		9'b110101101: rgb = 12'b010101010101;
		9'b110101110: rgb = 12'b010101010101;
		9'b110101111: rgb = 12'b000000000000;

		9'b110110000: rgb = 12'b000000000000;
		9'b110110001: rgb = 12'b100110011001;
		9'b110110010: rgb = 12'b100110011001;
		9'b110110011: rgb = 12'b010101010101;
		9'b110110100: rgb = 12'b110011001101;
		9'b110110101: rgb = 12'b110011001101;
		9'b110110110: rgb = 12'b010101010101;
		9'b110110111: rgb = 12'b010101010101;
		9'b110111000: rgb = 12'b010101010101;
		9'b110111001: rgb = 12'b010101010101;
		9'b110111010: rgb = 12'b010101010101;
		9'b110111011: rgb = 12'b100110011001;
		9'b110111100: rgb = 12'b100110011001;
		9'b110111101: rgb = 12'b010101010101;
		9'b110111110: rgb = 12'b010101010101;
		9'b110111111: rgb = 12'b000000000000;

		9'b111000000: rgb = 12'b000000000000;
		9'b111000001: rgb = 12'b010101010101;
		9'b111000010: rgb = 12'b010101010101;
		9'b111000011: rgb = 12'b010101010101;
		9'b111000100: rgb = 12'b110011001101;
		9'b111000101: rgb = 12'b110011001101;
		9'b111000110: rgb = 12'b010101010101;
		9'b111000111: rgb = 12'b010101010101;
		9'b111001000: rgb = 12'b010101010101;
		9'b111001001: rgb = 12'b010101010101;
		9'b111001010: rgb = 12'b010101010101;
		9'b111001011: rgb = 12'b100110011001;
		9'b111001100: rgb = 12'b100110011001;
		9'b111001101: rgb = 12'b010101010101;
		9'b111001110: rgb = 12'b010101010101;
		9'b111001111: rgb = 12'b000000000000;

		9'b111010000: rgb = 12'b000000000000;
		9'b111010001: rgb = 12'b010101010101;
		9'b111010010: rgb = 12'b010101010101;
		9'b111010011: rgb = 12'b010101010101;
		9'b111010100: rgb = 12'b010101010101;
		9'b111010101: rgb = 12'b010101010101;
		9'b111010110: rgb = 12'b010101010101;
		9'b111010111: rgb = 12'b010101010101;
		9'b111011000: rgb = 12'b010101010101;
		9'b111011001: rgb = 12'b010101010101;
		9'b111011010: rgb = 12'b010101010101;
		9'b111011011: rgb = 12'b010101010101;
		9'b111011100: rgb = 12'b010101010101;
		9'b111011101: rgb = 12'b010101010101;
		9'b111011110: rgb = 12'b000000000000;
		9'b111011111: rgb = 12'b000000000000;

		9'b111100000: rgb = 12'b000000000000;
		9'b111100001: rgb = 12'b000000000000;
		9'b111100010: rgb = 12'b010101010101;
		9'b111100011: rgb = 12'b010101010101;
		9'b111100100: rgb = 12'b010101010101;
		9'b111100101: rgb = 12'b010101010101;
		9'b111100110: rgb = 12'b010101010101;
		9'b111100111: rgb = 12'b010101010101;
		9'b111101000: rgb = 12'b010101010101;
		9'b111101001: rgb = 12'b010101010101;
		9'b111101010: rgb = 12'b010101010101;
		9'b111101011: rgb = 12'b010101010101;
		9'b111101100: rgb = 12'b010101010101;
		9'b111101101: rgb = 12'b000000000000;
		9'b111101110: rgb = 12'b000000000000;
		9'b111101111: rgb = 12'b000000000000;
		9'b111110000: rgb = 12'b011011011110;
		9'b111110001: rgb = 12'b000000000000;
		9'b111110010: rgb = 12'b000000000000;
		9'b111110011: rgb = 12'b000000000000;
		9'b111110100: rgb = 12'b000000000000;
		9'b111110101: rgb = 12'b000000000000;
		9'b111110110: rgb = 12'b000000000000;
		9'b111110111: rgb = 12'b000000000000;
		9'b111111000: rgb = 12'b000000000000;
		9'b111111001: rgb = 12'b000000000000;
		9'b111111010: rgb = 12'b000000000000;
		9'b111111011: rgb = 12'b000000000000;
		9'b111111100: rgb = 12'b000000000000;
		9'b111111101: rgb = 12'b000000000000;
		9'b111111110: rgb = 12'b000000000000;
		9'b111111111: rgb = 12'b011011011110;
		default: rgb = 12'b000000000000;
	endcase
endmodule